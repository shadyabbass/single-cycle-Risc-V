module data_memory(
    input         clk,
    input         wr_en,
    input  [31:0] addr,
    input  [31:0] write_data,
    output [31:0] read_data
    );

    // memory decleration
    reg [31:0] data_memory [2**31 -1:0];

initial
  begin
   data_memory [0]  =32'd0;
   data_memory [1]  =32'd1;
   data_memory [2]  =32'd2;
   data_memory [3]  =32'd3;
   data_memory [4]  =32'd4;
   data_memory [5]  =32'd5;
   data_memory [6]  =32'd6;
   data_memory [7]  =32'd7;
   data_memory [8]  =32'd8;
   data_memory [9]  =32'd9;
   data_memory [10] =32'd10;
   data_memory [11] =32'd11;
   data_memory [12] =32'd12;
   data_memory [13] =32'd13;
   data_memory [14] =32'd14;
   data_memory [15] =32'd15;
   data_memory [16] =32'd16;
   data_memory [17] =32'd17;
   data_memory [18] =32'd18;
   data_memory [19] =32'd19;
   data_memory [20] =32'd20;
   data_memory [21] =32'd21;
   data_memory [22] =32'd22;
   data_memory [23] =32'd23;
   data_memory [24] =32'd24;
   data_memory [25] =32'd25;
   data_memory [26] =32'd26;
   data_memory [27] =32'd27;
   data_memory [28] =32'd28;
   data_memory [29] =32'd29;
   data_memory [30] =32'd30;
   data_memory [31] =32'd31;
   data_memory [32] =32'd32;
   data_memory [33] =32'd33;
   data_memory [34] =32'd34;
   data_memory [35] =32'd35;
   data_memory [36] =32'd36;
   data_memory [37] =32'd37;
   data_memory [38] =32'd38;
   data_memory [39] =32'd39;
   data_memory [40] =32'd40;
   data_memory [41] =32'd41;
   data_memory [42] =32'd42;
   data_memory [43] =32'd43;
   data_memory [44] =32'd44;
   data_memory [45] =32'd45;
   data_memory [46] =32'd46;
   data_memory [47] =32'd47;
   data_memory [48] =32'd48;
   data_memory [49] =32'd49;
   data_memory [50] =32'd50;
   data_memory [51] =32'd51;
   data_memory [52] =32'd52;
   data_memory [53] =32'd53;
   data_memory [54] =32'd54;
   data_memory [55] =32'd55;
   data_memory [56] =32'd56;
   data_memory [57] =32'd57;
   data_memory [58] =32'd58;
   data_memory [59] =32'd59;
   data_memory [60] =32'd60;
   data_memory [61] =32'd61;
   data_memory [62] =32'd62;
   data_memory [63] =32'd63;
   data_memory [64] =32'd64;
   data_memory [65] =32'd65;
   data_memory [66] =32'd66;
   data_memory [67] =32'd67;
   data_memory [68] =32'd68;
   data_memory [69] =32'd69;
   data_memory [70] =32'd70;
   data_memory [71] =32'd71;
   data_memory [72] =32'd72;
   data_memory [73] =32'd73;
   data_memory [74] =32'd74;
   data_memory [75] =32'd75;
   data_memory [76] =32'd76;
   data_memory [77] =32'd77;
   data_memory [78] =32'd78;
   data_memory [79] =32'd79;
   data_memory [80] =32'd80;
   data_memory [81] =32'd81;
   data_memory [82] =32'd82;
   data_memory [83] =32'd83;
   data_memory [84] =32'd84;
   data_memory [85] =32'd85;
   data_memory [86] =32'd86;
   data_memory [87] =32'd87;
   data_memory [88] =32'd88;
   data_memory [89] =32'd89;
   data_memory [90] =32'd90;
   data_memory [91] =32'd91;
   data_memory [92] =32'd92;
   data_memory [93] =32'd93;
   data_memory [94] =32'd94;
   data_memory [95] =32'd95;
   data_memory [96] =32'd96;
   data_memory [97] =32'd97;
   data_memory [98] =32'd98;
   data_memory [99] =32'd99;
   data_memory [100]=32'd100;
   data_memory [101]=32'd101;
   data_memory [102]=32'd102;
   data_memory [103]=32'd103;
   data_memory [104]=32'd104;
   data_memory [105]=32'd105;
   data_memory [106]=32'd106;
   data_memory [107]=32'd107;
   data_memory [108]=32'd108;
   data_memory [109]=32'd109;
   data_memory [110]=32'd110;
   data_memory [111]=32'd111;
   data_memory [112]=32'd112;
   data_memory [113]=32'd113;
   data_memory [114]=32'd114;
   data_memory [115]=32'd115;
   data_memory [116]=32'd116;
   data_memory [117]=32'd117;
   data_memory [118]=32'd118;
   data_memory [119]=32'd119;
   data_memory [120]=32'd120;
   data_memory [121]=32'd121;
   data_memory [122]=32'd122;
   data_memory [123]=32'd123;
   data_memory [124]=32'd124;
   data_memory [125]=32'd125;
   data_memory [126]=32'd126;
   data_memory [127]=32'd127;
   data_memory [128]=32'd128;
   data_memory [129]=32'd129;
   data_memory [130]=32'd130;
   data_memory [131]=32'd131;
   data_memory [132]=32'd132;
   data_memory [133]=32'd133;
   data_memory [134]=32'd134;
   data_memory [135]=32'd135;
   data_memory [136]=32'd136;
   data_memory [137]=32'd137;
   data_memory [138]=32'd138;
   data_memory [139]=32'd139;
   data_memory [140]=32'd140;
   data_memory [141]=32'd141;
   data_memory [142]=32'd142;
   data_memory [143]=32'd143;
   data_memory [144]=32'd144;
   data_memory [145]=32'd145;
   data_memory [146]=32'd146;
   data_memory [147]=32'd147;
   data_memory [148]=32'd148;
   data_memory [149]=32'd149;
   data_memory [150]=32'd150;
   data_memory [151]=32'd151;
   data_memory [152]=32'd152;
   data_memory [153]=32'd153;
   data_memory [154]=32'd154;
   data_memory [155]=32'd155;
   data_memory [156]=32'd156;
   data_memory [157]=32'd157;
   data_memory [158]=32'd158;
   data_memory [159]=32'd159;
   data_memory [160]=32'd160;
   data_memory [161]=32'd161;
   data_memory [162]=32'd162;
   data_memory [163]=32'd163;
   data_memory [164]=32'd164;
   data_memory [165]=32'd165;
   data_memory [166]=32'd166;
   data_memory [167]=32'd167;
   data_memory [168]=32'd168;
   data_memory [169]=32'd169;
   data_memory [170]=32'd170;
   data_memory [171]=32'd171;
   data_memory [172]=32'd172;
   data_memory [173]=32'd173;
   data_memory [174]=32'd174;
   data_memory [175]=32'd175;
   data_memory [176]=32'd176;
   data_memory [177]=32'd177;
   data_memory [178]=32'd178;
   data_memory [179]=32'd179;
   data_memory [180]=32'd180;
   data_memory [181]=32'd181;
   data_memory [182]=32'd182;
   data_memory [183]=32'd183;
   data_memory [184]=32'd184;
   data_memory [185]=32'd185;
   data_memory [186]=32'd186;
   data_memory [187]=32'd187;
   data_memory [188]=32'd188;
   data_memory [189]=32'd189;
   data_memory [190]=32'd190;
   data_memory [191]=32'd191;
   data_memory [192]=32'd192;
   data_memory [193]=32'd193;
   data_memory [194]=32'd194;
   data_memory [195]=32'd195;
   data_memory [196]=32'd196;
   data_memory [197]=32'd197;
   data_memory [198]=32'd198;
   data_memory [199]=32'd199;
   data_memory [200]=32'd200;
   data_memory [201]=32'd201;
   data_memory [202]=32'd202;
   data_memory [203]=32'd203;
   data_memory [204]=32'd204;
   data_memory [205]=32'd205;
   data_memory [206]=32'd206;
   data_memory [207]=32'd207;
   data_memory [208]=32'd208;
   data_memory [209]=32'd209;
   data_memory [210]=32'd210;
   data_memory [211]=32'd211;
   data_memory [212]=32'd212;
   data_memory [213]=32'd213;
   data_memory [214]=32'd214;
   data_memory [215]=32'd215;
   data_memory [216]=32'd216;
   data_memory [217]=32'd217;
   data_memory [218]=32'd218;
   data_memory [219]=32'd219;
   data_memory [220]=32'd220;
   data_memory [221]=32'd221;
   data_memory [222]=32'd222;
   data_memory [223]=32'd223;
   data_memory [224]=32'd224;
   data_memory [225]=32'd225;
   data_memory [226]=32'd226;
   data_memory [227]=32'd227;
   data_memory [228]=32'd228;
   data_memory [229]=32'd229;
   data_memory [230]=32'd230;
   data_memory [231]=32'd231;
   data_memory [232]=32'd232;
   data_memory [233]=32'd233;
   data_memory [234]=32'd234;
   data_memory [235]=32'd235;
   data_memory [236]=32'd236;
   data_memory [237]=32'd237;
   data_memory [238]=32'd238;
   data_memory [239]=32'd239;
   data_memory [240]=32'd240;
   data_memory [241]=32'd241;
   data_memory [242]=32'd242;
   data_memory [243]=32'd243;
   data_memory [244]=32'd244;
   data_memory [245]=32'd245;
   data_memory [246]=32'd246;
   data_memory [247]=32'd247;
   data_memory [248]=32'd248;
   data_memory [249]=32'd249;
   data_memory [250]=32'd250;
   data_memory [251]=32'd251;
   data_memory [252]=32'd252;
   data_memory [253]=32'd253;
   data_memory [254]=32'd254;
   data_memory [255]=32'd255;
  end
    
    always@(posedge clk)
    begin
       if (wr_en) // case store instruction
          data_memory[addr[31:2]]<= write_data;
       else
          data_memory[addr[31:2]]<= data_memory[addr[31:2]];
    end
    
    assign read_data= data_memory[addr[31:2]]; 
endmodule
